library verilog;
use verilog.vl_types.all;
entity Frequency_Divider_vlg_vec_tst is
end Frequency_Divider_vlg_vec_tst;
