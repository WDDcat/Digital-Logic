library verilog;
use verilog.vl_types.all;
entity NameDispaly_vlg_vec_tst is
end NameDispaly_vlg_vec_tst;
