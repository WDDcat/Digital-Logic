library verilog;
use verilog.vl_types.all;
entity Selector_vlg_vec_tst is
end Selector_vlg_vec_tst;
