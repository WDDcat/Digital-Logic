library verilog;
use verilog.vl_types.all;
entity FlowLED_vlg_vec_tst is
end FlowLED_vlg_vec_tst;
