library verilog;
use verilog.vl_types.all;
entity Voter_vlg_vec_tst is
end Voter_vlg_vec_tst;
