library verilog;
use verilog.vl_types.all;
entity Chooser_vlg_vec_tst is
end Chooser_vlg_vec_tst;
