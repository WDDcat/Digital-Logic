library verilog;
use verilog.vl_types.all;
entity Scanner_vlg_vec_tst is
end Scanner_vlg_vec_tst;
