library verilog;
use verilog.vl_types.all;
entity Encoder_vlg_vec_tst is
end Encoder_vlg_vec_tst;
