library verilog;
use verilog.vl_types.all;
entity Shift_Reg_vlg_vec_tst is
end Shift_Reg_vlg_vec_tst;
