library verilog;
use verilog.vl_types.all;
entity Shift_Register_vlg_vec_tst is
end Shift_Register_vlg_vec_tst;
